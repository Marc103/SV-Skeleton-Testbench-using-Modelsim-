package golden_models_pkg;
    `include "ExampleModel.sv"
endpackage