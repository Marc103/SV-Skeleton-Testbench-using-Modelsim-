package generators_pkg;
    `include "ExampleGenerator.sv"
endpackage