package monitors_pkg;
    `include "ExampleMonitor.sv"
endpackage