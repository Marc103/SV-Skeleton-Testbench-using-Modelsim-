package scoreboards_pkg;
    `include "ExampleScoreboard.sv"
endpackage