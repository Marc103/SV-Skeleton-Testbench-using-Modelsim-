package utilities_pkg;
    `include "TriggerableQueue.sv"
    `include "TriggerableQueueBroadcaster.sv"
    `include "ExampleClass.sv"
endpackage