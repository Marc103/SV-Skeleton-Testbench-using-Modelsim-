package drivers_pkg;
    `include "ExampleDriver.sv"
endpackage